		
module C_NOT (a,c);
	input a;
	output c;
	
	assign c = !a;
endmodule 	